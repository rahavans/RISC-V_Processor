`timescale 1ns / 1ps

module RISCV_Processor();
endmodule